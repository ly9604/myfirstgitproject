`timescale 1ns / 1ps
module spi_ctrl #
  (
    
  )
